`timescale 1ns / 1ps

module Sumador_Serial();


endmodule
