`timescale 1ns / 1ps

module Main();
	//Este modulo se usara como principal para cargar y probar los proyectos. Este debe ser el modulo para la creacion del testbench.
	//Los modulos creados deben ser almacenados en nuevos archivos de Module Verilog.
	
	
endmodule
