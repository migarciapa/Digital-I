`timescale 1ns / 1ps

module Main(I,O);

	input I;
	output O;
	
	assign O = I;

endmodule
